class bridge_ahb_agent_config extends uvm_object;

	//Factory Registration
	`uvm_object_utils(bridge_ahb_agent_config)

        //Properties
	virtual ahb_if hvif;
	
	uvm_active_passive_enum is_active=UVM_ACTIVE;

	static int ahb_drv_data_count=0;
	static int ahb_mon_data_count=0;
		
		//------------------------------------------
		// Methods
		//------------------------------------------
		// Standard UVM Methods:
	extern function new(string name="bridge_ahb_agent_config");

endclass:bridge_ahb_agent_config

		//Constructor-new
function bridge_ahb_agent_config::new(string name="bridge_ahb_agent_config");
	super.new(name);
endfunction:new


